package uart_pkg;

    import uvm_pkg::*;
 
    `include "uvm_macros.svh"
 
    `include "typedefs.svh"
    `include "uart_seqit.svh"
 
    `include "uart_config.svh"
    `include "uart_driver.svh"
    `include "uart_monitor.svh"
    `include "uart_sequencer.svh"
    
    `include "uart_sequence.svh" 
 
    `include "uart_agent.svh"
 
 
 endpackage : uart_pkg