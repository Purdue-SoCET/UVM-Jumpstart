interface uart_if #(DATA_WIDTH = 8)
   (
   input reset,
   input clk
);
   // Bus Signals
endinterface