package uart_pkg;

endpackage : uart_pkg