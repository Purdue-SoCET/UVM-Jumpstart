package verif_pkg;

endpackage