`timescale 1ns/1ps
`include "uart_pkg.svh"
`include "uart_if.svh"
`include "verif_pkg.svh"
module top_tb;

   import uvm_pkg::*;
   import verif_pkg::*;

   initial
   begin
      // Initialize reset
   end

   // Clock Generation


   // Interface declarations

   // Connection of DUT
   initial
   begin
      // Register interfaces to uvm_config_db
      // Run UVM test class
   end

endmodule: top_tb