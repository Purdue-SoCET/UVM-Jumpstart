module top_tb;

   initial
   begin
      // Initialize reset
   end

   // Clock Generation


   // Interface declarations

   // Connection of DUT
   initial
   begin
      // Register interfaces to uvm_config_db
      // Run UVM test class
   end

endmodule: top_tb